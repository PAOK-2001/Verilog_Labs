module one_shot(

	input button, clock,
	output button_state
	
);


always @