module Full-Adder_tb();