module PinPlanner(
	
	//Switches
	input sw0, sw1, sw2, sw3, sw4, sw5, sw6, sw7, sw8, sw9,
	
	//Push_button
	input KEY0, KEY1,
	
	//Displays
	input[7:0] display_0, display_1, display_2, display_3, display_4, display_5,
	
	//LEDs
	input LEDR0, LEDR1, LEDR2, LEDR3, LEDR4, LEDR5, LEDR6, LEDR7, LEDR8, LEDR9,
	
	//miscelaneo
	input clk
	
);

endmodule
