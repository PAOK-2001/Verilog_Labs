module sum_tb();

endmodule
