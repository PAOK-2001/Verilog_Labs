module counter_tb();