module factorialSum_tb();