module Top_Level();

endmodule
